LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.display_types.ALL;
ENTITY encrypt IS

END encrypt;

ARCHITECTURE behavior OF encrypt IS
BEGIN

END behavior;