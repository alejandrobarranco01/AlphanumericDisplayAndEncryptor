LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY ascii_to_seven_segment IS
    PORT (
        ascii_in : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        seg_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END ascii_to_seven_segment;

ARCHITECTURE logic OF ascii_to_seven_segment IS
BEGIN
    PROCESS (ascii_in)
        VARIABLE H : STD_LOGIC := ascii_in(0); -- SW0
        VARIABLE G : STD_LOGIC := ascii_in(1); -- SW1
        VARIABLE F : STD_LOGIC := ascii_in(2); -- SW2
        VARIABLE E : STD_LOGIC := ascii_in(3); -- SW3
        VARIABLE D : STD_LOGIC := ascii_in(4); -- SW4
        VARIABLE C : STD_LOGIC := ascii_in(5); -- SW5
        VARIABLE B : STD_LOGIC := ascii_in(6); -- SW6
        VARIABLE A : STD_LOGIC := ascii_in(7); -- SW7
    BEGIN
        seg_out(0) <= NOT ((NOT A AND NOT B AND C AND D AND NOT E AND F AND H) OR (NOT A AND NOT B AND C AND D AND NOT E AND G) OR (NOT A AND NOT B AND C AND D AND E AND NOT F AND NOT G) OR (NOT A AND B AND NOT D AND NOT E AND F AND G) OR (NOT A AND B AND NOT D AND NOT F AND G AND H) OR (NOT A AND B AND NOT D AND F AND NOT G AND H) OR (NOT A AND B AND D AND NOT E AND NOT F AND NOT G) OR (NOT A AND B AND NOT E AND NOT F AND H) OR (NOT A AND B AND D AND E AND NOT F AND G AND NOT H) OR (NOT A AND NOT B AND C AND D AND NOT E AND NOT F AND NOT H));
        seg_out(1) <= NOT ((NOT A AND NOT B AND C AND D AND NOT E AND NOT F) OR (NOT A AND NOT B AND C AND D AND NOT E AND NOT G AND NOT H) OR (NOT A AND C AND D AND NOT F AND NOT G) OR (NOT A AND B AND NOT E AND NOT F AND NOT G AND H) OR (NOT A AND B AND NOT D AND NOT E AND F AND NOT G AND NOT H) OR (NOT A AND B AND E AND NOT F AND G AND NOT H) OR (NOT A AND B AND D AND NOT F AND NOT G) OR (NOT A AND B AND D AND NOT E AND F AND H) OR (NOT A AND NOT B AND C AND D AND NOT E AND G AND H));
        seg_out(2) <= NOT ((NOT A AND B AND NOT F AND NOT G AND H) OR (NOT A AND B AND NOT D AND NOT F AND G AND NOT H) OR (NOT A AND B AND NOT D AND NOT E AND F AND NOT G AND NOT H) OR (NOT A AND B AND NOT D AND F AND G AND H) OR (NOT A AND B AND NOT D AND E AND H) OR (NOT A AND B AND NOT D AND E AND G) OR (NOT A AND B AND D AND NOT E AND NOT F AND H) OR (NOT A AND B AND D AND NOT E AND NOT G AND H) OR (NOT A AND B AND D AND NOT E AND F AND G AND NOT H) OR (NOT A AND B AND E AND NOT F AND NOT G) OR (NOT A AND NOT B AND C AND D AND NOT F AND NOT G) OR (NOT A AND NOT B AND C AND D AND NOT E AND H) OR (NOT A AND NOT B AND C AND D AND NOT E AND F));
        seg_out(3) <= NOT ((NOT A AND C AND D AND NOT E AND F AND NOT G AND H) OR (NOT A AND NOT B AND C AND D AND NOT E AND G AND NOT H) OR (NOT A AND B AND NOT D AND F AND NOT G AND NOT H) OR (NOT A AND B AND NOT D AND F AND G AND H) OR (NOT A AND B AND NOT E AND G AND H) OR (NOT A AND B AND NOT E AND F AND NOT G) OR (NOT A AND B AND D AND E AND NOT F AND NOT G AND H) OR (NOT A AND B AND E AND NOT F AND G AND NOT H) OR (NOT A AND NOT B AND C AND D AND NOT E AND NOT F AND NOT H) OR (NOT A AND NOT B AND C AND D AND NOT E AND NOT F AND G) OR (NOT A AND NOT B AND C AND D AND E AND NOT F AND NOT G) OR (NOT A AND B AND NOT D AND NOT E AND NOT F AND G));
        seg_out(4) <= NOT ((NOT A AND C AND D AND NOT E AND G AND NOT H) OR (NOT A AND C AND D AND NOT F AND NOT G AND NOT H) OR (NOT A AND B AND NOT D AND NOT E AND H) OR (NOT A AND B AND NOT D AND G) OR (NOT A AND B AND NOT D AND F) OR (NOT A AND B AND NOT E AND F AND NOT G) OR (NOT A AND B AND E AND NOT F AND NOT H) OR (NOT A AND B AND D AND NOT E AND NOT H));
        seg_out(5) <= NOT ((NOT A AND C AND D AND NOT E AND F AND NOT G) OR (NOT A AND NOT B AND C AND D AND NOT E AND F AND NOT H) OR (NOT A AND C AND D AND E AND NOT F AND NOT G) OR (NOT A AND B AND NOT E AND H) OR (NOT A AND B AND NOT D AND NOT E AND G) OR (NOT A AND B AND NOT D AND NOT F AND G AND H) OR (NOT A AND B AND NOT D AND E AND NOT G AND NOT H) OR (NOT A AND B AND D AND NOT E AND NOT G) OR (NOT A AND B AND D AND NOT F AND NOT G) OR (NOT A AND C AND D AND NOT E AND NOT G AND NOT H));
        seg_out(6) <= NOT ((NOT A AND C AND D AND NOT E AND NOT F AND G) OR (NOT A AND NOT B AND C AND D AND NOT E AND F AND NOT G) OR (NOT A AND C AND D AND E AND NOT F AND NOT G) OR (NOT A AND B AND E AND NOT F AND NOT G AND NOT H) OR (NOT A AND B AND NOT D AND E AND G AND H) OR (NOT A AND B AND NOT D AND F AND G) OR (NOT A AND B AND D AND NOT E AND NOT F) OR (NOT A AND B AND D AND NOT F AND NOT G) OR (NOT A AND B AND D AND NOT F AND NOT H) OR (NOT A AND NOT B AND C AND D AND NOT E AND G AND NOT H) OR (NOT A AND B AND NOT D AND NOT E AND NOT G AND H) OR (NOT A AND B AND NOT D AND NOT E AND G AND NOT H) OR (NOT A AND B AND NOT E AND F AND NOT G AND NOT H));
    END PROCESS;
END logic;